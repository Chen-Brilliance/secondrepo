module moduleName (
    inout a
);
    
endmodule